magic
tech scmos
timestamp 1688669476
<< nwell >>
rect -28 -4 13 23
<< polysilicon >>
rect -9 11 -7 13
rect -9 -16 -7 1
rect -9 -23 -7 -21
<< ndiffusion >>
rect -19 -20 -17 -16
rect -13 -20 -9 -16
rect -19 -21 -9 -20
rect -7 -20 -4 -16
rect 0 -20 3 -16
rect -7 -21 3 -20
<< pdiffusion >>
rect -19 1 -17 11
rect -13 1 -9 11
rect -7 1 -4 11
rect 0 1 3 11
<< metal1 >>
rect -28 15 -25 19
rect -21 15 -17 19
rect -13 15 -9 19
rect -5 15 -1 19
rect 3 15 7 19
rect 11 15 13 19
rect -17 11 -13 15
rect -4 -8 0 1
rect -29 -12 -13 -8
rect -4 -12 14 -8
rect -4 -16 0 -12
rect -17 -26 -13 -20
rect -28 -30 -25 -26
rect -21 -30 -17 -26
rect -13 -30 -9 -26
rect -5 -30 -1 -26
rect 3 -30 7 -26
rect 11 -30 13 -26
<< ntransistor >>
rect -9 -21 -7 -16
<< ptransistor >>
rect -9 1 -7 11
<< polycontact >>
rect -13 -12 -9 -8
<< ndcontact >>
rect -17 -20 -13 -16
rect -4 -20 0 -16
<< pdcontact >>
rect -17 1 -13 11
rect -4 1 0 11
<< psubstratepcontact >>
rect -25 -30 -21 -26
rect -17 -30 -13 -26
rect -9 -30 -5 -26
rect -1 -30 3 -26
rect 7 -30 11 -26
<< nsubstratencontact >>
rect -25 15 -21 19
rect -17 15 -13 19
rect -9 15 -5 19
rect -1 15 3 19
rect 7 15 11 19
<< labels >>
rlabel metal1 5 17 5 17 1 vdd!
rlabel metal1 -11 -29 -11 -29 1 gnd!
rlabel metal1 -29 -12 -29 -8 3 vin
rlabel metal1 14 -12 14 -8 7 vout
<< end >>
